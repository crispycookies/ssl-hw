-- HPSPlatform_hmi.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HPSPlatform_hmi is
	port (
		leds_clk_clk                        : in  std_logic                     := '0';             --                     leds_clk.clk
		leds_external_connection_export     : out std_logic_vector(9 downto 0);                     --     leds_external_connection.export
		leds_reset_reset_n                  : in  std_logic                     := '0';             --                   leds_reset.reset_n
		leds_s1_address                     : in  std_logic_vector(1 downto 0)  := (others => '0'); --                      leds_s1.address
		leds_s1_write_n                     : in  std_logic                     := '0';             --                             .write_n
		leds_s1_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                             .writedata
		leds_s1_chipselect                  : in  std_logic                     := '0';             --                             .chipselect
		leds_s1_readdata                    : out std_logic_vector(31 downto 0);                    --                             .readdata
		seven_segment_clock_clk             : in  std_logic                     := '0';             --          seven_segment_clock.clk
		seven_segment_conduit_end_export    : out std_logic_vector(41 downto 0);                    --    seven_segment_conduit_end.export
		seven_segment_reset_reset           : in  std_logic                     := '0';             --          seven_segment_reset.reset
		seven_segment_s0_address            : in  std_logic_vector(7 downto 0)  := (others => '0'); --             seven_segment_s0.address
		seven_segment_s0_read               : in  std_logic                     := '0';             --                             .read
		seven_segment_s0_readdata           : out std_logic_vector(31 downto 0);                    --                             .readdata
		seven_segment_s0_write              : in  std_logic                     := '0';             --                             .write
		seven_segment_s0_writedata          : in  std_logic_vector(31 downto 0) := (others => '0'); --                             .writedata
		seven_segment_s0_waitrequest        : out std_logic;                                        --                             .waitrequest
		switches_clk_clk                    : in  std_logic                     := '0';             --                 switches_clk.clk
		switches_external_connection_export : in  std_logic_vector(9 downto 0)  := (others => '0'); -- switches_external_connection.export
		switches_reset_reset_n              : in  std_logic                     := '0';             --               switches_reset.reset_n
		switches_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  switches_s1.address
		switches_s1_readdata                : out std_logic_vector(31 downto 0)                     --                             .readdata
	);
end entity HPSPlatform_hmi;

architecture rtl of HPSPlatform_hmi is
	component HPSPlatform_hmi_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component HPSPlatform_hmi_leds;

	component seven_segment is
		port (
			avs_s0_address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_s0_read        : in  std_logic                     := 'X';             -- read
			avs_s0_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write       : in  std_logic                     := 'X';             -- write
			avs_s0_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_waitrequest : out std_logic;                                        -- waitrequest
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			seven_segment      : out std_logic_vector(41 downto 0)                     -- export
		);
	end component seven_segment;

	component HPSPlatform_hmi_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component HPSPlatform_hmi_switches;

begin

	leds : component HPSPlatform_hmi_leds
		port map (
			clk        => leds_clk_clk,                    --                 clk.clk
			reset_n    => leds_reset_reset_n,              --               reset.reset_n
			address    => leds_s1_address,                 --                  s1.address
			write_n    => leds_s1_write_n,                 --                    .write_n
			writedata  => leds_s1_writedata,               --                    .writedata
			chipselect => leds_s1_chipselect,              --                    .chipselect
			readdata   => leds_s1_readdata,                --                    .readdata
			out_port   => leds_external_connection_export  -- external_connection.export
		);

	seven_segment : component seven_segment
		port map (
			avs_s0_address     => seven_segment_s0_address,         --          s0.address
			avs_s0_read        => seven_segment_s0_read,            --            .read
			avs_s0_readdata    => seven_segment_s0_readdata,        --            .readdata
			avs_s0_write       => seven_segment_s0_write,           --            .write
			avs_s0_writedata   => seven_segment_s0_writedata,       --            .writedata
			avs_s0_waitrequest => seven_segment_s0_waitrequest,     --            .waitrequest
			clk                => seven_segment_clock_clk,          --       clock.clk
			reset              => seven_segment_reset_reset,        --       reset.reset
			seven_segment      => seven_segment_conduit_end_export  -- conduit_end.export
		);

	switches : component HPSPlatform_hmi_switches
		port map (
			clk      => switches_clk_clk,                    --                 clk.clk
			reset_n  => switches_reset_reset_n,              --               reset.reset_n
			address  => switches_s1_address,                 --                  s1.address
			readdata => switches_s1_readdata,                --                    .readdata
			in_port  => switches_external_connection_export  -- external_connection.export
		);

end architecture rtl; -- of HPSPlatform_hmi
